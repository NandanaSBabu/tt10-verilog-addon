`default_nettype none

module tt_um_addon (
    input  wire [7:0] ui_in,    // X input
    input  wire [7:0] uio_in,   // Y input
    output reg  [7:0] uo_out,   // Approximate Square Root Output
    output wire [7:0] uio_out,  // IOs: Output Path
    output wire [7:0] uio_oe,   // IOs: Enable Path
    input  wire        ena,      // Enable (ignored)
    input  wire        clk,      // Clock Signal
    input  wire        rst_n     // Active-low Reset
);

    assign uio_out = 8'b0;
    assign uio_oe  = 8'b0;

    // Define the LUT with an initial default value
    reg [7:0] sqrt_lut [0:65535];

    integer i;
    initial begin
        // Initialize entire LUT with zero to prevent 'x' values
        for (i = 0; i < 65536; i = i + 1) begin
            sqrt_lut[i] = 8'd0;
        end
        
        // Store values for specific (x, y) pairs
        sqrt_lut[(3  << 8) | 4]   = 8'd5;   // sqrt(3^2 + 4^2) = 5
        sqrt_lut[(5  << 8) | 12]  = 8'd13;  // sqrt(5^2 + 12^2) = 13
        sqrt_lut[(7  << 8) | 24]  = 8'd25;  // sqrt(7^2 + 24^2) = 25
        sqrt_lut[(8  << 8) | 15]  = 8'd17;  // sqrt(8^2 + 15^2) = 17
        sqrt_lut[(12 << 8) | 25]  = 8'd29;  // sqrt(12^2 + 25^2) = 29
        sqrt_lut[(9  << 8) | 40]  = 8'd41;  // sqrt(9^2 + 40^2) = 41
        sqrt_lut[(10 << 8) | 48]  = 8'd50;  // sqrt(10^2 + 48^2) = 50
        sqrt_lut[(11 << 8) | 60]  = 8'd61;  // sqrt(11^2 + 60^2) = 61
        sqrt_lut[(16 << 8) | 63]  = 8'd65;  // sqrt(16^2 + 63^2) = 65
        sqrt_lut[(13 << 8) | 84]  = 8'd85;  // sqrt(13^2 + 84^2) = 85
        sqrt_lut[(20 << 8) | 85]  = 8'd89;  // sqrt(20^2 + 85^2) = 89
        sqrt_lut[(48 << 8) | 55]  = 8'd97;  // sqrt(48^2 + 55^2) = 97
        sqrt_lut[(60 << 8) | 80]  = 8'd100; // sqrt(60^2 + 80^2) = 100
        sqrt_lut[(36 << 8) | 107] = 8'd113; // sqrt(36^2 + 107^2) = 113
        sqrt_lut[(35 << 8) | 115] = 8'd120; // sqrt(35^2 + 115^2) = 120
        sqrt_lut[(42 << 8) | 124] = 8'd130; // sqrt(42^2 + 124^2) = 130
        sqrt_lut[(70 << 8) | 120] = 8'd140; // sqrt(70^2 + 120^2) = 140
        sqrt_lut[(72 << 8) | 128] = 8'd145; // sqrt(72^2 + 128^2) = 145
        sqrt_lut[(80 << 8) | 137] = 8'd153; // sqrt(80^2 + 137^2) = 153
        sqrt_lut[(96 << 8) | 128] = 8'd160; // sqrt(96^2 + 128^2) = 160
    end

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            uo_out <= 8'd0;
        end else begin
            uo_out <= sqrt_lut[(ui_in << 8) | uio_in]; // Correct indexing using both X and Y
        end
    end

    wire _unused = &{ena, 1'b0};

endmodule
